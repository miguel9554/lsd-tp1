*******************************************************************************
** Circuito para simular el rise-time / fall-time de entrada de un flip-flop
** y en base a ello hacer una estimacion de su capacidad de entrada
*******************************************************************************

* Usar modelo del flip-flop lento, estando sus NMOS y PMOS dimensionados
* para que la excursion sea simetrica
.include ../caracteristicas_proceso/dig_0p25u_2p5V_stdcells_slow.inc

* Flip-flop cuya capacidad se va a analizar
* dff_x3ry1 RST D CLK QP VDD VSS
X1 0 2 4 5 4 0 dff_x3ry1


* Resistor que va entre la fuente cuadrada y el flip-flop
* Sirve para poder despejar Cin de la expresión de la
* constante de tiempo
R1 (1 2) r=1k

* Fuente de pulsos
vp 1 0 PULSE 2.5 0 0 0.1ps 0.1ps 3n 6n

* Alimentacion de 2.5V para el inversor
v1 4 0 dc 2.5

.end

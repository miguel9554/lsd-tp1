* Simulacion del rise-time y fall-time del inversor lento

.include inversor_clk.inc

X0 1 2 3 0 inversor_clk

** Fuentes
* Alimentacion
v1 3 0 dc 2.5

* Pulsos de entrada 
* Sintaxis: PULSE(V1 V2 DELAY RISE-TIME FALL-TIME DURACION_PULSO PERIODO)
vp 1 0 PULSE 0 2.5 0s 1ps 1ps 30n 60n
 
.end

**************************************************************************
*** Circuito para la simulacion del tiempo clock-to-Q la carga del FFD ***
**************************************************************************

** Cargar el inversor generador de la señal de clock
.include inversor_clk.inc

************ CIRCUITO ***************************************************

**** Descripcion de los nodos ****
* NODO 1: entrada de clk de flanco perfecto
* NODO 2: entrada de clk de FFD
* NODO 3: fuente de VCC=2.5V
* NODO 4: entrada D del FFD
* NODO 5: salida Q del FFD
*************************************************************************

** Fuente de alimentacion
v1 3 0 dc 2.5

** Senal de reloj
* Sintaxis: PULSE(V1 V2 DELAY RISE-TIME FALL-TIME DURACION_PULSO PERIODO)
vp_clk 1 0 PULSE 0 2.5 0s 30ps 30ps 50n 100n
X0 1 2 3 0 inversor_clk

** Flip-flop D
* NOTA: El reset se encuentra puesto a masa
X1 0 3 2 5 3 0 dff_x3ry1

.end

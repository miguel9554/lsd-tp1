
R1 1 2 10000.0
C1 2 0 1e-06

vp 1 0 PULSE 0 2.5 0 0 0 1 10

.end
